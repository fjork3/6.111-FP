/*
Parameterized module to generate Mel coefficient filter for 257-point FFT result (from 512-point transformation discarding negative frequencies).
To operate properly, requires that low, mid, and high are consecutive boundary points.
*/
module mel_filter(clock, coeffs);

   input clock;
   output [0:256] coeffs;

   // Parameters to determine start and end points for triangle filter.
   // 0 at low and high, maximum
   parameter low = 0;
   parameter mid = 9;
   parameter high = 16;
   

   // Implemented as 257-entry tables, with 2 entries for each index.
   // Assumes fixed placements of bin edges, as determined by Mel scale.
   // Based on low, mid, and high, assigns entry 0, 1023, or table entry.

   wire [0:256] ascending [9:0];
   wire [0:256] descending [9:0];

   for (i=0; i<257; i=i+1) begin
      assign ascending[i] = 10'h2AA;
   end  
   
   


/*
   if ((i > low) && (i <= mid)) 
      coeffs[i] <= ascending[i];
   else if ((i > mid) && (i < high))
      coeffs[i] <= descending[i];
   else
      coeffs[i] <= 10'b0;
*/

   // Values generated with python (create_coeffs.py)
   assign ascending[0] = 1023;
   assign ascending[1] = 341;
   assign ascending[2] = 682;
   assign ascending[3] = 1023;
   assign ascending[4] = 341;
   assign ascending[5] = 682;
   assign ascending[6] = 1023;
   assign ascending[7] = 256;
   assign ascending[8] = 512;
   assign ascending[9] = 767;
   assign ascending[10] = 1023;
   assign ascending[11] = 256;
   assign ascending[12] = 512;
   assign ascending[13] = 767;
   assign ascending[14] = 1023;
   assign ascending[15] = 256;
   assign ascending[16] = 512;
   assign ascending[17] = 767;
   assign ascending[18] = 1023;
   assign ascending[19] = 171;
   assign ascending[20] = 341;
   assign ascending[21] = 512;
   assign ascending[22] = 682;
   assign ascending[23] = 853;
   assign ascending[24] = 1023;
   assign ascending[25] = 171;
   assign ascending[26] = 341;
   assign ascending[27] = 512;
   assign ascending[28] = 682;
   assign ascending[29] = 853;
   assign ascending[30] = 1023;
   assign ascending[31] = 171;
   assign ascending[32] = 341;
   assign ascending[33] = 512;
   assign ascending[34] = 682;
   assign ascending[35] = 853;
   assign ascending[36] = 1023;
   assign ascending[37] = 128;
   assign ascending[38] = 256;
   assign ascending[39] = 384;
   assign ascending[40] = 512;
   assign ascending[41] = 639;
   assign ascending[42] = 767;
   assign ascending[43] = 895;
   assign ascending[44] = 1023;
   assign ascending[45] = 128;
   assign ascending[46] = 256;
   assign ascending[47] = 384;
   assign ascending[48] = 512;
   assign ascending[49] = 639;
   assign ascending[50] = 767;
   assign ascending[51] = 895;
   assign ascending[52] = 1023;
   assign ascending[53] = 102;
   assign ascending[54] = 205;
   assign ascending[55] = 307;
   assign ascending[56] = 409;
   assign ascending[57] = 512;
   assign ascending[58] = 614;
   assign ascending[59] = 716;
   assign ascending[60] = 818;
   assign ascending[61] = 921;
   assign ascending[62] = 1023;
   assign ascending[63] = 102;
   assign ascending[64] = 205;
   assign ascending[65] = 307;
   assign ascending[66] = 409;
   assign ascending[67] = 512;
   assign ascending[68] = 614;
   assign ascending[69] = 716;
   assign ascending[70] = 818;
   assign ascending[71] = 921;
   assign ascending[72] = 1023;
   assign ascending[73] = 79;
   assign ascending[74] = 157;
   assign ascending[75] = 236;
   assign ascending[76] = 315;
   assign ascending[77] = 393;
   assign ascending[78] = 472;
   assign ascending[79] = 551;
   assign ascending[80] = 630;
   assign ascending[81] = 708;
   assign ascending[82] = 787;
   assign ascending[83] = 866;
   assign ascending[84] = 944;
   assign ascending[85] = 1023;
   assign ascending[86] = 79;
   assign ascending[87] = 157;
   assign ascending[88] = 236;
   assign ascending[89] = 315;
   assign ascending[90] = 393;
   assign ascending[91] = 472;
   assign ascending[92] = 551;
   assign ascending[93] = 630;
   assign ascending[94] = 708;
   assign ascending[95] = 787;
   assign ascending[96] = 866;
   assign ascending[97] = 944;
   assign ascending[98] = 1023;
   assign ascending[99] = 64;
   assign ascending[100] = 128;
   assign ascending[101] = 192;
   assign ascending[102] = 256;
   assign ascending[103] = 320;
   assign ascending[104] = 384;
   assign ascending[105] = 448;
   assign ascending[106] = 512;
   assign ascending[107] = 575;
   assign ascending[108] = 639;
   assign ascending[109] = 703;
   assign ascending[110] = 767;
   assign ascending[111] = 831;
   assign ascending[112] = 895;
   assign ascending[113] = 959;
   assign ascending[114] = 1023;
   assign ascending[115] = 60;
   assign ascending[116] = 120;
   assign ascending[117] = 181;
   assign ascending[118] = 241;
   assign ascending[119] = 301;
   assign ascending[120] = 361;
   assign ascending[121] = 421;
   assign ascending[122] = 481;
   assign ascending[123] = 542;
   assign ascending[124] = 602;
   assign ascending[125] = 662;
   assign ascending[126] = 722;
   assign ascending[127] = 782;
   assign ascending[128] = 842;
   assign ascending[129] = 903;
   assign ascending[130] = 963;
   assign ascending[131] = 1023;
   assign ascending[132] = 54;
   assign ascending[133] = 108;
   assign ascending[134] = 162;
   assign ascending[135] = 215;
   assign ascending[136] = 269;
   assign ascending[137] = 323;
   assign ascending[138] = 377;
   assign ascending[139] = 431;
   assign ascending[140] = 485;
   assign ascending[141] = 538;
   assign ascending[142] = 592;
   assign ascending[143] = 646;
   assign ascending[144] = 700;
   assign ascending[145] = 754;
   assign ascending[146] = 808;
   assign ascending[147] = 861;
   assign ascending[148] = 915;
   assign ascending[149] = 969;
   assign ascending[150] = 1023;
   assign ascending[151] = 44;
   assign ascending[152] = 89;
   assign ascending[153] = 133;
   assign ascending[154] = 178;
   assign ascending[155] = 222;
   assign ascending[156] = 267;
   assign ascending[157] = 311;
   assign ascending[158] = 356;
   assign ascending[159] = 400;
   assign ascending[160] = 445;
   assign ascending[161] = 489;
   assign ascending[162] = 534;
   assign ascending[163] = 578;
   assign ascending[164] = 623;
   assign ascending[165] = 667;
   assign ascending[166] = 712;
   assign ascending[167] = 756;
   assign ascending[168] = 801;
   assign ascending[169] = 845;
   assign ascending[170] = 890;
   assign ascending[171] = 934;
   assign ascending[172] = 979;
   assign ascending[173] = 1023;
   assign ascending[174] = 43;
   assign ascending[175] = 85;
   assign ascending[176] = 128;
   assign ascending[177] = 171;
   assign ascending[178] = 213;
   assign ascending[179] = 256;
   assign ascending[180] = 298;
   assign ascending[181] = 341;
   assign ascending[182] = 384;
   assign ascending[183] = 426;
   assign ascending[184] = 469;
   assign ascending[185] = 512;
   assign ascending[186] = 554;
   assign ascending[187] = 597;
   assign ascending[188] = 639;
   assign ascending[189] = 682;
   assign ascending[190] = 725;
   assign ascending[191] = 767;
   assign ascending[192] = 810;
   assign ascending[193] = 853;
   assign ascending[194] = 895;
   assign ascending[195] = 938;
   assign ascending[196] = 980;
   assign ascending[197] = 1023;
   assign ascending[198] = 37;
   assign ascending[199] = 73;
   assign ascending[200] = 110;
   assign ascending[201] = 146;
   assign ascending[202] = 183;
   assign ascending[203] = 219;
   assign ascending[204] = 256;
   assign ascending[205] = 292;
   assign ascending[206] = 329;
   assign ascending[207] = 365;
   assign ascending[208] = 402;
   assign ascending[209] = 438;
   assign ascending[210] = 475;
   assign ascending[211] = 512;
   assign ascending[212] = 548;
   assign ascending[213] = 585;
   assign ascending[214] = 621;
   assign ascending[215] = 658;
   assign ascending[216] = 694;
   assign ascending[217] = 731;
   assign ascending[218] = 767;
   assign ascending[219] = 804;
   assign ascending[220] = 840;
   assign ascending[221] = 877;
   assign ascending[222] = 913;
   assign ascending[223] = 950;
   assign ascending[224] = 986;
   assign ascending[225] = 1023;
   assign ascending[226] = 33;
   assign ascending[227] = 66;
   assign ascending[228] = 99;
   assign ascending[229] = 132;
   assign ascending[230] = 165;
   assign ascending[231] = 198;
   assign ascending[232] = 231;
   assign ascending[233] = 264;
   assign ascending[234] = 297;
   assign ascending[235] = 330;
   assign ascending[236] = 363;
   assign ascending[237] = 396;
   assign ascending[238] = 429;
   assign ascending[239] = 462;
   assign ascending[240] = 495;
   assign ascending[241] = 528;
   assign ascending[242] = 561;
   assign ascending[243] = 594;
   assign ascending[244] = 627;
   assign ascending[245] = 660;
   assign ascending[246] = 693;
   assign ascending[247] = 726;
   assign ascending[248] = 759;
   assign ascending[249] = 792;
   assign ascending[250] = 825;
   assign ascending[251] = 858;
   assign ascending[252] = 891;
   assign ascending[253] = 924;
   assign ascending[254] = 957;
   assign ascending[255] = 990;
   assign ascending[256] = 1023;
   
   assign descending[0] = 1023;
   assign descending[1] = 682;
   assign descending[2] = 341;
   assign descending[3] = 1023;
   assign descending[4] = 682;
   assign descending[5] = 341;
   assign descending[6] = 1023;
   assign descending[7] = 767;
   assign descending[8] = 511;
   assign descending[9] = 256;
   assign descending[10] = 1023;
   assign descending[11] = 767;
   assign descending[12] = 511;
   assign descending[13] = 256;
   assign descending[14] = 1023;
   assign descending[15] = 767;
   assign descending[16] = 511;
   assign descending[17] = 256;
   assign descending[18] = 1023;
   assign descending[19] = 852;
   assign descending[20] = 682;
   assign descending[21] = 511;
   assign descending[22] = 341;
   assign descending[23] = 170;
   assign descending[24] = 1023;
   assign descending[25] = 852;
   assign descending[26] = 682;
   assign descending[27] = 511;
   assign descending[28] = 341;
   assign descending[29] = 170;
   assign descending[30] = 1023;
   assign descending[31] = 852;
   assign descending[32] = 682;
   assign descending[33] = 511;
   assign descending[34] = 341;
   assign descending[35] = 170;
   assign descending[36] = 1023;
   assign descending[37] = 895;
   assign descending[38] = 767;
   assign descending[39] = 639;
   assign descending[40] = 511;
   assign descending[41] = 384;
   assign descending[42] = 256;
   assign descending[43] = 128;
   assign descending[44] = 1023;
   assign descending[45] = 895;
   assign descending[46] = 767;
   assign descending[47] = 639;
   assign descending[48] = 511;
   assign descending[49] = 384;
   assign descending[50] = 256;
   assign descending[51] = 128;
   assign descending[52] = 1023;
   assign descending[53] = 921;
   assign descending[54] = 818;
   assign descending[55] = 716;
   assign descending[56] = 614;
   assign descending[57] = 511;
   assign descending[58] = 409;
   assign descending[59] = 307;
   assign descending[60] = 205;
   assign descending[61] = 102;
   assign descending[62] = 1023;
   assign descending[63] = 921;
   assign descending[64] = 818;
   assign descending[65] = 716;
   assign descending[66] = 614;
   assign descending[67] = 511;
   assign descending[68] = 409;
   assign descending[69] = 307;
   assign descending[70] = 205;
   assign descending[71] = 102;
   assign descending[72] = 1023;
   assign descending[73] = 944;
   assign descending[74] = 866;
   assign descending[75] = 787;
   assign descending[76] = 708;
   assign descending[77] = 630;
   assign descending[78] = 551;
   assign descending[79] = 472;
   assign descending[80] = 393;
   assign descending[81] = 315;
   assign descending[82] = 236;
   assign descending[83] = 157;
   assign descending[84] = 79;
   assign descending[85] = 1023;
   assign descending[86] = 944;
   assign descending[87] = 866;
   assign descending[88] = 787;
   assign descending[89] = 708;
   assign descending[90] = 630;
   assign descending[91] = 551;
   assign descending[92] = 472;
   assign descending[93] = 393;
   assign descending[94] = 315;
   assign descending[95] = 236;
   assign descending[96] = 157;
   assign descending[97] = 79;
   assign descending[98] = 1023;
   assign descending[99] = 959;
   assign descending[100] = 895;
   assign descending[101] = 831;
   assign descending[102] = 767;
   assign descending[103] = 703;
   assign descending[104] = 639;
   assign descending[105] = 575;
   assign descending[106] = 511;
   assign descending[107] = 448;
   assign descending[108] = 384;
   assign descending[109] = 320;
   assign descending[110] = 256;
   assign descending[111] = 192;
   assign descending[112] = 128;
   assign descending[113] = 64;
   assign descending[114] = 1023;
   assign descending[115] = 963;
   assign descending[116] = 903;
   assign descending[117] = 842;
   assign descending[118] = 782;
   assign descending[119] = 722;
   assign descending[120] = 662;
   assign descending[121] = 602;
   assign descending[122] = 542;
   assign descending[123] = 481;
   assign descending[124] = 421;
   assign descending[125] = 361;
   assign descending[126] = 301;
   assign descending[127] = 241;
   assign descending[128] = 181;
   assign descending[129] = 120;
   assign descending[130] = 60;
   assign descending[131] = 1023;
   assign descending[132] = 969;
   assign descending[133] = 915;
   assign descending[134] = 861;
   assign descending[135] = 808;
   assign descending[136] = 754;
   assign descending[137] = 700;
   assign descending[138] = 646;
   assign descending[139] = 592;
   assign descending[140] = 538;
   assign descending[141] = 485;
   assign descending[142] = 431;
   assign descending[143] = 377;
   assign descending[144] = 323;
   assign descending[145] = 269;
   assign descending[146] = 215;
   assign descending[147] = 162;
   assign descending[148] = 108;
   assign descending[149] = 54;
   assign descending[150] = 1023;
   assign descending[151] = 979;
   assign descending[152] = 934;
   assign descending[153] = 890;
   assign descending[154] = 845;
   assign descending[155] = 801;
   assign descending[156] = 756;
   assign descending[157] = 712;
   assign descending[158] = 667;
   assign descending[159] = 623;
   assign descending[160] = 578;
   assign descending[161] = 534;
   assign descending[162] = 489;
   assign descending[163] = 445;
   assign descending[164] = 400;
   assign descending[165] = 356;
   assign descending[166] = 311;
   assign descending[167] = 267;
   assign descending[168] = 222;
   assign descending[169] = 178;
   assign descending[170] = 133;
   assign descending[171] = 89;
   assign descending[172] = 44;
   assign descending[173] = 1023;
   assign descending[174] = 980;
   assign descending[175] = 938;
   assign descending[176] = 895;
   assign descending[177] = 852;
   assign descending[178] = 810;
   assign descending[179] = 767;
   assign descending[180] = 725;
   assign descending[181] = 682;
   assign descending[182] = 639;
   assign descending[183] = 597;
   assign descending[184] = 554;
   assign descending[185] = 511;
   assign descending[186] = 469;
   assign descending[187] = 426;
   assign descending[188] = 384;
   assign descending[189] = 341;
   assign descending[190] = 298;
   assign descending[191] = 256;
   assign descending[192] = 213;
   assign descending[193] = 170;
   assign descending[194] = 128;
   assign descending[195] = 85;
   assign descending[196] = 43;
   assign descending[197] = 1023;
   assign descending[198] = 986;
   assign descending[199] = 950;
   assign descending[200] = 913;
   assign descending[201] = 877;
   assign descending[202] = 840;
   assign descending[203] = 804;
   assign descending[204] = 767;
   assign descending[205] = 731;
   assign descending[206] = 694;
   assign descending[207] = 658;
   assign descending[208] = 621;
   assign descending[209] = 585;
   assign descending[210] = 548;
   assign descending[211] = 511;
   assign descending[212] = 475;
   assign descending[213] = 438;
   assign descending[214] = 402;
   assign descending[215] = 365;
   assign descending[216] = 329;
   assign descending[217] = 292;
   assign descending[218] = 256;
   assign descending[219] = 219;
   assign descending[220] = 183;
   assign descending[221] = 146;
   assign descending[222] = 110;
   assign descending[223] = 73;
   assign descending[224] = 37;
   assign descending[225] = 1023;
   assign descending[226] = 990;
   assign descending[227] = 957;
   assign descending[228] = 924;
   assign descending[229] = 891;
   assign descending[230] = 858;
   assign descending[231] = 825;
   assign descending[232] = 792;
   assign descending[233] = 759;
   assign descending[234] = 726;
   assign descending[235] = 693;
   assign descending[236] = 660;
   assign descending[237] = 627;
   assign descending[238] = 594;
   assign descending[239] = 561;
   assign descending[240] = 528;
   assign descending[241] = 495;
   assign descending[242] = 462;
   assign descending[243] = 429;
   assign descending[244] = 396;
   assign descending[245] = 363;
   assign descending[246] = 330;
   assign descending[247] = 297;
   assign descending[248] = 264;
   assign descending[249] = 231;
   assign descending[250] = 198;
   assign descending[251] = 165;
   assign descending[252] = 132;
   assign descending[253] = 99;
   assign descending[254] = 66;
   assign descending[255] = 33;
   assign descending[256] = 0;


endmodule //mel_filter
