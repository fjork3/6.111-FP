/*
Main voice control module.
*/
module voice_control_main (
   // Inputs


   // Outputs

)






endmodule
