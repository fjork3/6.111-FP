/*///////////////////////////////////////////////////////////////////////////////

Main video filter module.

*////////////////////////////////////////////////////////////////////////////////
module video_filter_main (clk, vclk, fvh, dv, ntsc_addr, ntsc_data, ntsc_we, sw)

   // Inputs
   input 	 clk;

   ///////////////////////////////////////////////////////////////////////////////
   // Outputs

   ///////////////////////////////////////////////////////////////////////////////
   // NTSC video interface

   input 	 vclk;	// video clock from camera
   input [2:0] 	 fvh;
   input 	 dv;
   input [7:0] 	 din;
   output [18:0] ntsc_addr;
   output [35:0] ntsc_data;
   output 	 ntsc_we;	// write enable for NTSC data
   input 	 sw;		// switch which determines mode (for debugging)



   ///////////////////////////////////////////////////////////////////////////////
   // NTSC conversion


   // instantiate zbt_6111

   // instantiate ntsc2zbt


endmodule
