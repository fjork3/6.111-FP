
module filter_mult(clock, filter, score, fft_data, start, done);

   input clock;
   


endmodule
